module BirdROM(
    input clka,
    input ena,
    input [10:0] addra,
    output [11:0] douta
);
endmodule
