module PillarMainROM(
    input clka,
    input ena,
    input [5:0] addra,
    output [11:0] douta
);
endmodule
