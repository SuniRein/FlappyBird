module BackgroundInitROM(
    input clka,
    input ena,
    input [18:0] addra,
    output [11:0] douta
);
endmodule
