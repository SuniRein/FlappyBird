module SongROM(
    input clka,
    input ena,
    input [7:0] addra,
    output douta
);
endmodule
