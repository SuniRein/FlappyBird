module Display
#(
    parameter WIDTH  = 640,
    parameter HEIGHT = 480
)
(
    input clk,
    input rstn

);



endmodule
